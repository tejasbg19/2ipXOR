** sch_path: /home/tejas/Desktop/Github/2ipXOR/Schematic Simulation/threshold/nmoss_threshold.sch
**.subckt nmoss_threshold
VCC VCC GND 5
R1 VCC Vo 1k m=1
Vinn Vinn GND 0
XM1 Vo Vinn GND GND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.dc Vinn -10 10 1
.save all
.end

**** end user architecture code
**.ends
.GLOBAL GND
.end
